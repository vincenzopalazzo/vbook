module markdown

pub struct MDDocument {

}