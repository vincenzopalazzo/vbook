module markdown

struct Scanner { }

pub fn (instance &Scanner) scan() ([]&Token) {
	return []&Token{}
}